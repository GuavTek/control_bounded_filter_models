package Coefficients;
	localparam real Lfr[0:2] = {0.9742006659182473, 0.9510703751817556, 0.9742006659182456};
	localparam real Lfi[0:2] = {0.04199890731649758, 2.800111352637899e-15, -0.04199890731649972};
	localparam real Lbr[0:2] = {0.9742006659182415, 0.9510703751817727, 0.9742006659182332};
	localparam real Lbi[0:2] = {0.04199890731648781, 1.3469880457339309e-14, -0.04199890731650077};
	localparam real Wfr[0:2] = {-3.857664364797836e-07, -0.00016579813393585724, -3.8576643643676786e-07};
	localparam real Wfi[0:2] = {-0.00028862319171261714, -4.2666350772185406e-19, 0.0002886231917126176};
	localparam real Wbr[0:2] = {3.764739916262334e-07, 0.0001664613896363954, 3.7647399140998926e-07};
	localparam real Wbi[0:2] = {0.00028919709182248813, -1.7457011560855188e-18, -0.0002891970918224965};
localparam real Ffr[0:2][0:59] = '{
	'{24.47889595448819, -2.272267731204669, -0.040102784734557945, 23.222083180140405, -2.2769723024217097, -0.028353204258878825, 21.970648454207193, -2.2759136180947985, -0.017112456216094328, 20.727367720601254, -2.269377624713338, -0.0063828312989029495, 19.494860622183385, -2.2576495162179024, 0.0038347342121347744, 18.275591821494338, -2.241013078119799, 0.013540594128003375, 17.07187263307436, -2.2197500672915154, 0.022736328058933594, 15.88586294808396, -2.1941396271809435, 0.03142467730520509, 14.719573432177938, -2.164457738128388, 0.03960948107780217, 13.574867977857242, -2.130976702395828, 0.047295613187656696, 12.453466392828155, -2.093964663452801, 0.05448891933425236, 11.35694730623316, -2.053685159002434, 0.061196155116478676, 10.286751274980158, -2.010396707174585, 0.06742492488082559, 9.244184072784474, -1.9643524252606341, 0.07318362151431658, 8.230420144949168, -1.9157996803161794, 0.07848136728200217, 7.246506212340827, -1.8649797709135778, 0.08332795580138978, 6.293365008469275, -1.8121276392859118, 0.08773379523888195, 5.371799134047177, -1.7574716130674015, 0.09170985280614213, 4.482495013888543, -1.7012331758024892, 0.09526760062731959, 3.626026941500821, -1.643626765366605, 0.09841896304124464},
	'{-48.53773741100753, 4.38418921246969, -0.4000303614506594, -46.16280412996046, 4.1696724791713535, -0.38045702594897196, -43.9040754433234, 3.965651969150541, -0.3618414064098237, -41.75586550388969, 3.7716141061402726, -0.3441366421504851, -39.7127666708233, 3.5870704429676312, -0.32729816536385153, -37.76963589712543, 3.4115564319966114, -0.31128358892889857, -35.92158178315739, 3.244630255732749, -0.29605259971053094, -34.16395226362962, 3.0858717146458217, -0.28156685708022877, -32.49232289706181, 2.934881169410969, -0.267789896402041, -30.902485728235327, 2.79127853490556, -0.2546870372409726, -29.390438695601624, 2.654702323429412, -0.24222529606270157, -27.952375556982222, 2.524808734739889, -0.2303733032048654, -26.58467630820042, 2.4012707906112407, -0.21910122391091172, -25.283898070525705, 2.2837775117396233, -0.20838068322773265, -24.04676642399215, 2.1720331349218602, -0.19818469457803026, -22.87016716477426, 2.0657563685373383, -0.1884875918276089, -21.751138465871325, 1.9646796844589076, -0.17926496467658962, -20.686863421366557, 1.8685486446103063, -0.17049359721190827, -19.674662955492828, 1.7771212604748852, -0.16215140946641673, -18.711989078655154, 1.6901673839433236, -0.15421740183747543},
	'{24.478895954487243, -2.272267731204316, -0.040102784734594214, 23.222083180139634, -2.276972302421374, -0.028353204258913717, 21.970648454206586, -2.2759136180944792, -0.01711245621612786, 20.72736772060081, -2.269377624713035, -0.0063828312989351425, 19.494860622183086, -2.2576495162176142, 0.00383473421210391, 18.275591821494185, -2.2410130781195257, 0.013540594127973815, 17.071872633074342, -2.2197500672912556, 0.02273632805890531, 15.885862948084071, -2.194139627180697, 0.031424677305178034, 14.719573432178166, -2.1644577381281542, 0.03960948107777634, 13.574867977857583, -2.130976702395607, 0.04729561318763204, 12.453466392828602, -2.0939646634525912, 0.054488919334228836, 11.356947306233714, -2.053685159002236, 0.06119615511645627, 10.286751274980801, -2.0103967071743973, 0.06742492488080427, 9.244184072785211, -1.964352425260457, 0.07318362151429629, 8.230420144949985, -1.9157996803160113, 0.07848136728198285, 7.246506212341726, -1.8649797709134197, 0.08332795580137142, 6.293365008470247, -1.8121276392857624, 0.08773379523886449, 5.371799134048218, -1.7574716130672607, 0.09170985280612556, 4.48249501388965, -1.7012331758023564, 0.09526760062730381, 3.626026941501988, -1.6436267653664802, 0.09841896304122968}};
localparam real Ffi[0:2][0:59] = '{
	'{14.88785303278273, 1.5078384078030567, -0.25512462155163523, 15.53184322103267, 1.3735044191377144, -0.250226849346944, 16.106434128046555, 1.2424385710739754, -0.2449619668622122, 16.613642081222935, 1.1147985981960642, -0.2393608157043881, 17.0555479746673, 0.9907261562008656, -0.23345353799408927, 17.434289038940616, 0.8703472683287374, -0.22726953752805373, 17.752050878612227, 0.7537727878229712, -0.2208374446449697, 18.01105978379418, 0.6410988745062265, -0.21418508469794892, 18.21357532086482, 0.532407483621978, -0.20733945003290594, 18.361883206655083, 0.4277668651502592, -0.20032667536853896, 18.45828846947218, 0.32723207186960535, -0.19317201647047388, 18.50510889947241, 0.23084547450080217, -0.18589983200941088, 18.504668790068543, 0.13863728233268557, -0.1785335684907954, 18.45929297126714, 0.05062606779558099, -0.17109574814160233, 18.371301135077985, -0.03318070648618121, -0.16360795963826427, 18.243002452421177, -0.11278615956505078, -0.15609085155857394, 18.076690480277456, -0.1882034643003765, -0.14856412843953326, 17.874638357183933, -0.2594553210175803, -0.14104654932259494, 17.63909428457012, -0.32657343389995275, -0.1335559286675281, 17.372277290857927, -0.3895979912508222, -0.12610913951622393},
	'{-5.335218159580759e-12, 2.062032721767128e-13, 4.145517467174695e-15, -5.210079006264908e-12, 2.083900414187609e-13, 2.8225492963305246e-15, -5.084412787128856e-12, 2.0986914212199206e-13, 1.6191209806795043e-15, -4.958570677109478e-12, 2.1070459083646544e-13, 5.26701768616897e-16, -4.832870747280426e-12, 2.1095583373572814e-13, -4.626904698568923e-16, -4.7076003636205596e-12, 2.1067804060788454e-13, -1.3565225072926954e-15, -4.583018430294915e-12, 2.0992238101889646e-13, -2.1617770812030373e-15, -4.459357486921215e-12, 2.0873628368887898e-13, -2.884982385106513e-15, -4.3368256687401e-12, 2.0716368006299148e-13, -3.53223983243293e-15, -4.215608538084155e-12, 2.0524523300265333e-13, -4.10925019170101e-15, -4.095870795047472e-12, 2.0301855147006393e-13, -4.621338185884941e-15, -3.977757874792357e-12, 2.0051839202919914e-13, -5.07347564369261e-15, -3.861397438491254e-12, 1.977768479394373e-13, -5.470303285570866e-15, -3.746900764488543e-12, 1.9482352657357398e-13, -5.816151222615678e-15, -3.6343640458771442e-12, 1.91685715850083e-13, -6.1150582421833366e-15, -3.523869600317511e-12, 1.8838854032992223e-13, -6.370789949858608e-15, -3.4154869975803698e-12, 1.849551075908479e-13, -6.586855833524051e-15, -3.3092741099682555e-12, 1.814066454569601e-13, -6.766525311579006e-15, -3.2052780904634177e-12, 1.7776263062794427e-13, -6.912842823865428e-15, -3.1035362831599035e-12, 1.7404090922108468e-13, -7.028642020559351e-15},
	'{-14.887853032777343, -1.5078384078032647, 0.255124621551631, -15.53184322102741, -1.3735044191379244, 0.2502268493469411, -16.10643412804142, -1.242438571074187, 0.24496196686221042, -16.613642081217932, -1.1147985981962767, 0.23936081570438741, -17.055547974662417, -0.9907261562010785, 0.2334535379940895, -17.43428903893586, -0.8703472683289506, 0.22726953752805487, -17.752050878607598, -0.7537727878231837, 0.22083744464497163, -18.011059783789676, -0.6410988745064388, 0.2141850846979516, -18.213575320860436, -0.5324074836221889, 0.20733945003290918, -18.361883206650823, -0.427766865150469, 0.20032667536854276, -18.45828846946804, -0.32723207186981385, 0.19317201647047816, -18.50510889946839, -0.23084547450100912, 0.18589983200941562, -18.504668790064642, -0.1386372823328904, 0.17853356849080051, -18.459292971263356, -0.050626067795783936, 0.17109574814160775, -18.371301135074315, 0.03318070648598048, 0.16360795963826993, -18.243002452417628, 0.11278615956485194, 0.15609085155857982, -18.076690480274017, 0.18820346430017998, 0.1485641284395393, -17.874638357180604, 0.25945532101738633, 0.1410465493226011, -17.6390942845669, 0.3265734338997609, 0.13355592866753435, -17.37227729085482, 0.389597991250633, 0.12610913951623026}};
localparam real Fbr[0:2][0:59] = '{
	'{-24.430836501043682, -2.756372996107157, -0.05947710737410642, -23.176540121016707, -2.7359868347330485, -0.07093974034516513, -21.927608707916793, -2.7099559257516583, -0.08166641626485872, -20.686812767029128, -2.678621059083147, -0.09166726091124705, -19.45676681499454, -2.6423191543341895, -0.1009536656035808, -18.23993069763487, -2.6013826325471654, -0.10953819730134347, -17.038611218756774, -2.5561388297692313, -0.11743451026741322, -15.854964060686438, -2.5069094518097756, -0.1246572594330535, -14.690995977524839, -2.454010069485724, -0.13122201559153643, -13.548567242385776, -2.397749653590263, -0.13714518253652427, -12.429394330182808, -2.338430148761597, -0.14244391625090075, -11.335052817865575, -2.276346085374372, -0.1471360462415651, -10.266980484367497, -2.211784228527113, -0.15123999910579167, -9.226480592913859, -2.1450232631545054, -0.15477472440512788, -8.214725338749359, -2.0763335142533093, -0.15775962291346074, -7.232759445775281, -2.0059767011751113, -0.1602144772968389, -6.281503896036457, -1.934205724907828, -0.16215938527389662, -5.361759776465069, -1.8612644872407387, -0.16361469529729875, -4.4742122277701295, -1.7873877406846934, -0.1646009447885129, -3.6194344808563947, -1.712800967999918, -0.165138800950423},
	'{48.34434162659983, 5.333510489909506, 0.5943941974630557, 45.97887112872609, 5.072543822674155, 0.5653107123870571, 43.7291422148319, 4.824346156556692, 0.5376502713242336, 41.589491692637274, 4.588292709123117, 0.5113432452649207, 39.55453346773576, 4.363789268309515, 0.48632341212077346, 37.61914498529943, 4.1502706966253236, 0.46252779002538386, 35.77845433518623, 3.947199508545364, 0.439896478791438, 34.0278279879895, 3.7540645175095486, 0.41837250912531376, 32.362859131158, 3.570379549124387, 0.39790169921955176, 30.779356575825297, 3.3956822173270593, 0.378432518362204, 29.273334206423726, 3.22953276043132, 0.3599159572197244, 27.841000946524836, 3.071512934125242, 0.3423054044668702, 26.478751215647467, 2.9212249586341614, 0.3255565294530547, 25.183155853010657, 2.7782905173985504, 0.30962717060979256, 23.950953485383902, 2.642349804746201, 0.2944772293183262, 22.779042317305258, 2.5130606201614536, 0.28006856897026944, 21.664472323000986, 2.390097506871492, 0.2663649189671763, 20.604437820351677, 2.2731509325812893, 0.25333178341737483, 19.59627040821138, 2.1619265102948835, 0.24093635430023033, 18.637432249301067, 2.0561442572615753, 0.22914742887924858},
	'{-24.430836501038648, -2.756372996105259, -0.059477107373856246, -23.176540121012568, -2.7359868347312624, -0.07093974034492644, -21.927608707913507, -2.7099559257499792, -0.08166641626463125, -20.68681276702664, -2.6786210590815696, -0.09166726091103052, -19.45676681499281, -2.6423191543327094, -0.1009536656033749, -18.239930697633845, -2.601382632545778, -0.1095381973011479, -17.038611218756422, -2.5561388297679324, -0.11743451026722765, -15.85496406068671, -2.5069094518085597, -0.12465725943287757, -14.690995977525706, -2.454010069484588, -0.13122201559136984, -13.5485672423872, -2.397749653589202, -0.13714518253636665, -12.429394330184753, -2.338430148760608, -0.14244391625075173, -11.335052817868004, -2.2763460853734503, -0.14713604624142432, -10.266980484370386, -2.2117842285262554, -0.15123999910565877, -9.22648059291718, -2.1450232631537087, -0.1547747244050025, -8.21472533875308, -2.0763335142525703, -0.15775962291334256, -7.232759445779377, -2.0059767011744256, -0.16021447729672753, -6.281503896040905, -1.9342057249071942, -0.16215938527379176, -5.361759776469845, -1.8612644872401534, -0.16361469529720005, -4.4742122277752125, -1.7873877406841538, -0.16460094478842, -3.6194344808617602, -1.712800967999422, -0.1651388009503356}};
localparam real Fbi[0:2][0:59] = '{
	'{-14.857459565257917, 1.2078034798415764, 0.3094628780810575, -15.500215440199211, 1.060878300366859, 0.2989809683834839, -16.07370956417772, 0.9185998891845217, 0.28828806691625836, -16.57995416699435, 0.7810854359985733, 0.277420526518524, -17.021025922455813, 0.6484347942924246, 0.26641333687876745, -17.399057734409574, 0.5207310911407759, 0.2553001065518516, -17.716230790040864, 0.39804134767460664, 0.2441130492157375, -17.9747668865973, 0.2804171081680428, 0.23288297399282573, -18.17692103673926, 0.1678950757947888, 0.22163927965957514, -18.324974356781638, 0.0604977531816181, 0.2104099525672858, -18.421227241195535, -0.0417659140331883, 0.19922156809662117, -18.467992825877367, -0.13889989234773514, 0.18809929546858548, -18.467590741868065, -0.23092041588102374, 0.17706690573523406, -18.42234116041656, -0.31785534374339053, 0.16614678277435768, -18.334559129530007, -0.3997435207614187, 0.15535993711372673, -18.206549201438044, -0.47663414294551887, 0.14472602241218224, -18.040600349719735, -0.5485861290085821, 0.13426335442689677, -17.838981174199617, -0.6156674991650951, 0.12398893229848267, -17.60393539111327, -0.677954762361948, 0.11391846198826694, -17.33767760547266, -0.7355323130150957, 0.10406638170497245},
	'{2.7409497429793943e-11, 1.6506795635511478e-12, 3.567140000577867e-14, 2.6719553506597034e-11, 1.6417541805285213e-12, 4.1932430571118504e-14, 2.6031505675876043e-11, 1.6297503233375404e-12, 4.74953601926643e-14, 2.534682018783765e-11, 1.614990617482893e-12, 5.2413514920424135e-14, 2.4666815267093014e-11, 1.5977734867796678e-12, 5.673667368634965e-14, 2.399267208796986e-11, 1.578374749312177e-12, 6.051128775431455e-14, 2.3325445030178042e-11, 1.55704911515491e-12, 6.37806871870674e-14, 2.266607125897658e-11, 1.5340315916482023e-12, 6.658527507528065e-14, 2.2015379671392776e-11, 1.5095388016895406e-12, 6.896271023198378e-14, 2.137409924759511e-11, 1.4837702201883495e-12, 7.094807901614424e-14, 2.0742866844212912e-11, 1.4569093335365836e-12, 7.25740569118191e-14, 2.01222344642194e-11, 1.429124726668536e-12, 7.387106045402565e-14, 1.9512676035943104e-11, 1.4005711020200314e-12, 7.486739005915553e-14, 1.891459373183919e-11, 1.3713902344487381e-12, 7.558936428628008e-14, 1.8328323855829707e-11, 1.3417118659428986e-12, 7.606144602596219e-14, 1.775414232630441e-11, 1.3116545437245543e-12, 7.630636108510639e-14, 1.71922697802557e-11, 1.2813264051446103e-12, 7.634520960985556e-14, 1.66428763224962e-11, 1.2508259125701404e-12, 7.619757076349315e-14, 1.6106085942471125e-11, 1.2202425412785262e-12, 7.588160105265172e-14, 1.558198061982419e-11, 1.1896574231977525e-12, 7.541412667279032e-14},
	'{14.8574595652302, -1.2078034798432453, -0.3094628780810935, 15.500215440172191, -1.0608783003685187, -0.29898096838352617, 16.073709564151397, -0.9185998891861696, -0.2882880669163062, 16.57995416696872, -0.7810854360002063, -0.2774205265185766, 17.02102592243087, -0.6484347942940405, -0.2664133368788244, 17.399057734385313, -0.5207310911423725, -0.25530010655191215, 17.716230790017278, -0.3980413476761828, -0.24411304921580126, 17.97476688657438, -0.280417108169596, -0.232882973992892, 18.176921036717, -0.16789507579631824, -0.2216392796596436, 18.32497435676003, -0.06049775318312278, -0.21040995256735598, 18.42122724117457, 0.041765914031709706, -0.19922156809669261, 18.46799282585703, 0.13889989234628353, -0.18809929546865783, 18.467590741848355, 0.23092041587959888, -0.177066905735307, 18.42234116039746, 0.31785534374199287, -0.16614678277443093, 18.334559129511504, 0.39974352076004915, -0.15535993711379997, 18.206549201420124, 0.47663414294417683, -0.14472602241225518, 18.040600349702398, 0.5485861290072683, -0.13426335442696924, 17.838981174182848, 0.615667499163809, -0.1239889322985545, 17.603935391097053, 0.6779547623606895, -0.11391846198833788, 17.33767760545699, 0.7355323130138647, -0.1040663817050424}};
	localparam real hf[0:1199] = {0.09036497, -0.0025117926, -0.009208244, 0.085569896, -0.008494271, -0.00834019, 0.07845638, -0.013158934, -0.006855863, 0.06969149, -0.016434716, -0.0050614374, 0.059936076, -0.01837167, -0.0031910879, 0.049796417, -0.019103622, -0.0014145782, 0.039793197, -0.018816262, 0.00015411813, 0.030344823, -0.017720906, 0.0014477256, 0.021762133, -0.01603382, 0.0024365978, 0.014251728, -0.013960793, 0.0031200734, 0.00792538, -0.011686433, 0.0035185567, 0.0028133253, -0.009367564, 0.0036665378, -0.0011204077, -0.007130022, 0.0036066615, -0.003962103, -0.005068188, 0.0033848952, -0.005833038, -0.0032465511, 0.0030467694, -0.0068755466, -0.0017027154, 0.0026346256, -0.0072409683, -0.0004513, 0.002185764, -0.007079774, 0.0005117207, 0.0017313665, -0.0065339375, 0.0012046016, 0.0012960604, -0.0057314746, 0.0016556147, 0.00089798385, -0.004782968, 0.0018992391, 0.0005492241, -0.003779821, 0.001972879, 0.00025650932, -0.0027939335, 0.0019141743, 2.205085e-05, -0.0018785027, 0.0017589165, -0.00015555069, -0.0010696395, 0.0015395507, -0.00028040342, -0.00038852476, 0.0012842063, -0.00035847822, 0.00015613581, 0.0010161905, -0.000396854, 0.000565563, 0.0007538644, -0.0004030763, 0.00084842165, 0.00051081745, -0.0003846385, 0.0010185246, 0.0002962626, -0.00034858685, 0.0010928051, 0.0001155782, -0.00030124193, 0.0010896028, -2.9068606e-05, -0.00024802543, 0.0010272873, -0.00013806968, -0.00019337657, 0.0009232092, -0.00021373798, -0.00014074247, 0.0007929628, -0.00025971574, -9.262507e-05, 0.00064992433, -0.00028045053, -5.066916e-05, 0.00050502596, -0.00028075196, -1.5776592e-05, 0.0003667219, -0.00026543438, 1.1765581e-05, 0.00024110163, -0.00023904513, 3.2153504e-05, 0.00013210971, -0.00020567249, 4.5939545e-05, 4.1833468e-05, -0.00016882573, 5.3915883e-05, -2.9173532e-05, -0.00013137597, 5.7012578e-05, -8.1558894e-05, -9.5547155e-05, 5.6212357e-05, -0.00011685057, -6.2945364e-05, 5.2482843e-05, -0.00013716304, -3.4615852e-05, 4.6725843e-05, -0.00014494038, -1.1117832e-05, 3.9742452e-05, -0.0001427421, 7.391287e-06, 3.2212123e-05, -0.00013307319, 2.1069243e-05, 2.4683577e-05, -0.00011825778, 3.0305251e-05, 1.7575183e-05, -0.00010035267, 3.5643305e-05, 1.1182553e-05, -8.1096485e-05, 3.7715057e-05, 5.691199e-06, -6.188855e-05, 3.7183774e-05, 1.1923481e-06, -4.379175e-05, 3.4699857e-05, -2.2997494e-06, -2.7553384e-05, 3.0867643e-05, -4.830316e-06, -1.3638718e-05, 2.6222673e-05, -6.487387e-06, -2.2722415e-06, 2.1218233e-05, -7.386724e-06, 6.5174827e-06, 1.6219634e-05, -7.658765e-06, 1.2852708e-05, 1.1504807e-05, -7.4378595e-06, 1.6963733e-05, 7.269602e-06, -6.8538516e-06, 1.915029e-05, 3.6364115e-06, -6.025907e-06, 1.9748253e-05, 6.648429e-07, -5.0584126e-06, 1.910227e-05, -1.6366539e-06, -4.0386717e-06, 1.7544417e-05, -3.29907e-06, -3.036102e-06, 1.537864e-05, -4.3817104e-06, -2.102623e-06, 1.2870485e-05, -4.9621394e-06, -1.2739252e-06, 1.0241401e-05, -5.1274983e-06, -5.7134537e-07, 7.666878e-06, -4.9673586e-06, -4.0933723e-09, 5.2775918e-06, -4.5681404e-06, 4.2837235e-07, 3.16277e-06, -4.009039e-06, 7.339921e-07, 1.3750837e-06, -3.3593205e-06, 9.258993e-07, -6.359334e-08, -2.676821e-06, 1.02045e-06, -1.1560729e-06, -2.0074363e-06, 1.0355419e-06, -1.9238194e-06, -1.3854044e-06, 9.892484e-07, -2.4013098e-06, -8.341688e-07, 8.9876687e-07, -2.6310133e-06, -3.676398e-07, 7.7966735e-07, -2.6591165e-06, 8.312268e-09, 6.4541064e-07, -2.5320603e-06, 2.9427056e-07, 5.0709895e-07, -2.2938889e-06, 4.957026e-07, 3.734177e-07, -1.9843594e-06, 6.2149206e-07, 2.5072586e-07, -1.6377461e-06, 6.8262983e-07, 1.432551e-07, -1.2822309e-06, 6.910985e-07, 5.3379903e-08, -9.3978184e-07, 6.589672e-07, -1.8072758e-08, -6.264063e-07, 5.97698e-07, -7.150114e-08, -3.5267666e-07, 5.1764965e-07, -1.0821479e-07, -1.2443446e-07, 4.277629e-07, -1.3014446e-07, 5.640928e-08, 3.3539862e-07, -1.3958638e-07, 1.910447e-07, 2.4630316e-07, -1.3898715e-07, 2.8295824e-07, 1.6467209e-07, -1.3077126e-07, 3.3719118e-07, 9.32852e-08, -1.1721109e-07, 3.5968802e-07, 3.368847e-08, -1.0033626e-07, 3.567494e-07, -1.3598448e-08, -8.187813e-08, 3.3459582e-07, -4.8866845e-08, -6.324415e-08, 2.9903916e-07, -7.30096e-08, -4.551648e-08, 2.552557e-07, -8.7328075e-08, -2.946897e-08, 2.076485e-07, -9.336221e-08, -1.5597422e-08, 1.5978559e-07, -9.274775e-08, -4.158099e-09, 1.1439974e-07, -8.710208e-08, 4.789537e-09, 7.3434734e-08, -7.793836e-08, 1.1339283e-08, 3.812472e-08, -6.660583e-08, 1.5696466e-08, 9.094313e-09, -5.4253537e-08, 1.8139922e-08, -1.35311655e-08, -4.1813852e-08, 1.8988922e-08, -3.0013776e-08, -3.0002017e-08, 1.8575733e-08, -4.08961e-08, -1.9327915e-08, 1.7223961e-08, -4.690415e-08, -1.0116509e-08, 1.5232557e-08, -4.8863175e-08, -2.5337308e-09, 1.2864989e-08, -4.7627942e-08, 3.384918e-09, 1.0342998e-08, -4.4028017e-08, 7.705285e-09, 7.844139e-09, -3.8827427e-08, 1.05667635e-08, 5.502401e-09, -3.2697635e-08, 1.2156995e-08, 3.4110983e-09, -2.6202096e-08, 1.2689909e-08, 1.627343e-09, -1.979051e-08, 1.2387518e-08, 1.7748072e-10, -1.3800811e-08, 1.1465601e-08, -9.370555e-10, -8.466915e-09, 1.0123142e-08, -1.7338936e-09, -3.9304298e-09, 8.5352205e-09, -2.2441988e-09, -2.5472774e-10, 6.84893e-09, -2.5077114e-09, 2.5599607e-09, 5.1818296e-09, -2.5684856e-09, 4.5615254e-09, 3.6224153e-09, -2.4714037e-09, 5.8318466e-09, 2.232099e-09, -2.2594735e-09, 6.4741275e-09, 1.0482302e-09, -1.9718722e-09, 6.602058e-09, 8.7739704e-11, -1.6426741e-09, 6.3309704e-09, -6.489429e-10, -1.3001609e-09, 5.77101e-09, -1.1739845e-09, -9.666239e-10, 5.0222204e-09, -1.5084695e-09, -6.585453e-10, 4.1713655e-09, -1.6790994e-09, -3.8706144e-10, 3.2902467e-09, -1.7153653e-09, -1.5861411e-10, 2.4352584e-09, -1.6472363e-09, 2.429134e-11, 1.6479078e-09, -1.5033739e-09, 1.6228845e-10, 9.560427e-10, -1.3098419e-09, 2.5836688e-10, 3.7554979e-10, -1.0892715e-09, 3.1714453e-10, -8.768451e-11, -8.604138e-10, 3.44222e-10, -4.357213e-10, -6.3801825e-10, 3.4563594e-10, -6.7656175e-10, -4.329611e-10, 3.2741826e-10, -8.2228596e-10, -2.525611e-10, 2.9526048e-10, -8.874075e-10, -1.01017764e-10, 2.5427718e-10, -8.874836e-10, 2.008026e-11, 2.0885768e-10, -8.379982e-10, 1.1122219e-10, 1.6259383e-10, -7.535152e-10, 1.7445302e-10, 1.1826932e-10, -6.470841e-10, 2.1288897e-10, 7.789677e-11, -5.298726e-10, 2.3028836e-10, 4.278894e-11, -4.1099088e-10, 2.3068897e-10, 1.36521e-11, -2.974732e-10, 2.181161e-10, -9.308972e-12, -1.9437936e-10, 1.9636077e-10, -2.6283024e-11, -1.0498246e-10, 1.6882395e-10, -3.7748082e-11, -3.101161e-11, 1.3841953e-10, -4.437588e-11, 2.7076966e-11, 1.07527605e-10, -4.694825e-11, 6.982229e-11, 7.798881e-11, -4.6287238e-11, 9.849156e-11, 5.1129923e-11, -4.319966e-11, 1.1483604e-10, 2.7812206e-11, -3.8435675e-11, 1.2087802e-10, 8.49416e-12, -3.2660413e-11, 1.1873334e-10, -6.6981737e-12, -2.6437066e-11, 1.1047113e-10, -1.789908e-11, -2.0219751e-11, 9.800927e-11, -2.5433688e-11, -1.43541064e-11, 8.3043426e-11, -2.975438e-11, -9.083842e-12, 6.7005304e-11, -3.1385228e-11, -4.5614003e-12, 5.1045546e-11, -3.0875687e-11, -8.6117685e-13, 3.6036434e-11, -2.8763854e-11, 2.0060468e-12, 2.2589486e-11, -2.5549151e-11, 4.0785582e-12, 1.1083396e-11, -2.1673644e-11, 5.4298926e-12, 1.6983405e-12, -1.7511029e-11, 6.156334e-12, -5.546812e-12, -1.3362047e-11, 6.366126e-12, -1.0757145e-11, -9.455064e-12, 6.1705775e-12, -1.4126313e-11, -5.950565e-12, 5.6771224e-12, -1.590464e-11, -2.9483482e-12, 4.9842435e-12, -1.6371656e-11, -4.964109e-13, 4.1781058e-12, -1.581353e-11, 1.399398e-12, 3.33068e-12, -1.4505517e-11, 2.7656677e-12, 2.4991042e-12, -1.2699198e-11, 3.652218e-12, 1.7260272e-12, -1.0614062e-11, 4.1237846e-12, 1.040676e-12, -8.432901e-12, 4.2528567e-12, 4.6042114e-13, -6.3003426e-12, 4.1137814e-12, -7.36975e-15, -4.3238624e-12, 3.778172e-12, -3.633617e-13, -2.576632e-12, 3.311561e-12, -6.1430255e-13, -1.1016023e-12, 2.7711906e-12, -7.711978e-13, 8.369866e-14, 2.2047897e-12, -8.4768233e-13, 9.820906e-13, 1.6501753e-12, -8.586334e-13, 1.6117382e-12, 1.1355021e-12, -8.190441e-13, 2.0014836e-12, 6.799909e-13, -7.4315884e-13, 2.1866933e-12, 2.949831e-13, -6.4385644e-13, 2.205731e-12, -1.4816282e-14, -5.3225637e-13, 2.0971016e-12, -2.50021e-13, -4.1751685e-13, 1.8972688e-12, -4.1526293e-13, -3.0679075e-13, 1.639105e-12, -5.179766e-13, -2.0530364e-13, 1.3509112e-12, -5.6731697e-13, -1.1652105e-13, 1.0559265e-12, -5.732385e-13, -4.237409e-14, 7.722352e-13, -5.4574926e-13, 1.6482958e-14, 5.1298505e-13, -4.943395e-13, 6.040517e-14, 2.8682886e-13, -4.2757478e-13, 9.049681e-14, 9.8511504e-14, -3.5283853e-13, 1.0837127e-13, -5.0464227e-14, -2.76201e-13, 1.1593981e-13, -1.6114962e-13, -2.0239314e-13, 1.1523389e-13, -2.364832e-13, -1.3486147e-13, 1.0826318e-13, -2.8067723e-13, -7.588145e-14, 9.690856e-14, -2.986794e-13, -2.6709351e-14, 8.284776e-14, -2.9572137e-13, 1.22452275e-14, 6.751009e-14, -2.769592e-13, 4.1240594e-14, 5.2055826e-14, -2.4720344e-13, 6.102953e-14, 3.737544e-14, -2.1073295e-13, 7.2699496e-14, 2.4104196e-14, -1.7118251e-13, 7.753227e-14, 1.2647414e-14, -1.3149341e-13, 7.6886095e-14, 3.2126153e-15, -9.391428e-14, 7.210166e-14, -4.1549698e-15, -6.004055e-14, 6.443142e-14, -9.536281e-15, -3.088089e-14, 5.499072e-14, -1.3103869e-14, -6.9406384e-15, 4.4728154e-14, -1.509045e-14, 1.1686564e-14, 3.441232e-14, -1.5761579e-14, 2.5225974e-14, 2.4631779e-14, -1.5393021e-14, 3.4133236e-14, 1.5805064e-14, -1.4252915e-14, 3.9014083e-14, 8.1978026e-15, -1.2588622e-14, 4.0554792e-14, 1.9442976e-15, -1.0617867e-14, 3.9464685e-14, -2.9287005e-15, -8.523638e-15, 3.6431053e-14, -6.4778767e-15, -6.4522472e-15, 3.2086025e-14, -8.820321e-15, -4.51389e-15, 2.6984422e-14, -1.0112606e-14, -2.7850964e-15, 2.159119e-14, -1.053265e-14, -1.3124761e-15, 1.6276843e-14, -1.0264695e-14, -1.1723878e-16, 1.1319271e-14, -9.487522e-15, 7.9994067e-16, 6.910272e-15, -8.365769e-15, 1.4540708e-15, 3.1653545e-15, -7.0441064e-15, 1.8712705e-15, 1.3544979e-16, -5.643916e-15, 2.0846665e-15, -2.180554e-15, -4.262062e-15, 2.1308744e-15, -3.823357e-15, -2.9713185e-15, 2.0471247e-15, -4.8615486e-15, -1.8220469e-15, 1.8690373e-15, -5.381139e-15, -8.44718e-16, 1.6290167e-15, -5.476608e-15, -5.2948728e-17, 1.3552095e-15, -5.243616e-15, 5.5324513e-16, 1.0709456e-15, -4.77338e-15, 9.842112e-16, 7.945839e-16, -4.1486424e-15, 1.2576151e-15, 5.396705e-16, -3.4410677e-15, 1.3957121e-15, 3.1532874e-16, -2.7098803e-15, 1.4230113e-15, 1.2680276e-16, -2.0015213e-15, 1.3643713e-15, -2.3911259e-17, -1.3500983e-15, 1.243529e-15, -1.3740334e-16, -7.784197e-16, 1.0820415e-15, -2.1620091e-16, -2.994108e-16, 8.98602e-16, -2.641664e-16, 8.2253894e-17, 7.08678e-16, -2.8596364e-16, 3.6844713e-16, 5.2441594e-16, -2.866069e-16, 5.659254e-16, 3.5475397e-16, -2.7109732e-16, 6.8478887e-16, 2.0568692e-16, -2.441469e-16, 7.371213e-16, 8.0632435e-17, -2.0998436e-16, 7.358432e-16, -1.9146106e-17, -1.7223414e-16, 6.937914e-16, -9.409717e-17, -1.3385789e-16, 6.230221e-16, -1.4594842e-16, -9.7146996e-17, 5.343241e-16, -1.7730566e-16, -6.37543e-17, 4.3691796e-16, -1.9129831e-16, -3.4753815e-17, 3.3831483e-16, -1.9128e-16, -1.07186345e-17, 2.443042e-16, -1.8058791e-16, 8.191798e-18, 1.5904068e-16, -1.6236055e-16, 2.2142091e-17, 8.520121e-17, -1.3940967e-16, 3.1534554e-17, 2.4187628e-17, -1.1414125e-16, 3.693014e-17, -2.3648035e-17, -8.85177e-17, 3.8979358e-17, -5.877322e-17, -6.405402e-17, 3.8364624e-17, -8.225363e-17, -4.1839705e-17, 3.575458e-17, -9.555126e-17, -2.2579241e-17, 3.1770042e-17, -1.00348437e-16, -6.644488e-18, 2.6960733e-17, -9.840144e-17, 5.8669046e-18, 2.1791517e-17, -9.142484e-17, 1.5071644e-17, 1.6636663e-17, -8.100571e-17, 2.124324e-17, 1.1780518e-17, -6.8545427e-17, 2.47594e-17, 7.423046e-18, -5.5225592e-17, 2.6056133e-17, 3.688762e-18, -4.1994454e-17, 2.5589525e-17, 6.3773904e-19, -2.9569517e-17, 2.38055e-17, -1.7223943e-18, -1.8452424e-17, 2.1117347e-17, -3.4243954e-18, -8.952369e-18, 1.7890414e-17, -4.529961e-18, -1.2146473e-18, 1.4433135e-17, -5.1193935e-18, 4.7484224e-18, 1.0993361e-17, -5.2826864e-18, 9.026524e-18, 7.758946e-18, -5.1121937e-18, 1.178205e-17, 4.86155e-18, -4.696912e-18, 1.3223719e-17, 2.3826712e-18, -4.118312e-18, 1.3583899e-17, 3.610363e-19, -3.4475817e-18, 1.31000015e-17, -1.1993739e-18, -2.7441022e-18, 1.2000025e-17, -2.3212744e-18, -2.0549429e-18, 1.0492073e-17, -3.0464508e-18, -1.4151657e-18, 8.757471e-18, -3.428886e-18, -8.4872753e-19, 6.94702e-18, -3.5288422e-18, -3.6978636e-19, 5.179849e-18, -3.4080017e-18, 1.5755416e-20, 3.544303e-18, -3.125685e-18, 3.086148e-19, 2.1003448e-18, -2.736102e-18, 5.1451203e-19, 8.829621e-19, -2.2865427e-18, 6.426599e-19, -9.3835756e-20, -1.8163844e-18, 7.044178e-19, -8.328061e-19, -1.3567788e-18, 7.1214657e-19, -1.3493264e-18, -9.308701e-19, 6.7827973e-19, -1.6675306e-18, -5.544108e-19, 6.1461246e-19, -1.8168768e-18, -2.3664195e-19, 5.317948e-19, -1.8292355e-18, 1.8672093e-20, 4.3901003e-19, -1.7365352e-18, 2.1214996e-19, 3.4381106e-19, -1.5689669e-18, 3.477149e-19, 2.520872e-19, -1.3537122e-18, 4.3158893e-19, 1.6813144e-19, -1.1141423e-18, 4.713982e-19, 9.4780856e-20, -8.694209e-19, 4.754127e-19, 3.3604972e-20, -6.3443605e-19, 4.5193163e-19, -1.4880066e-20, -4.199873e-19, 4.0881287e-19, -5.098947e-20, -2.331562e-19, 3.5313953e-19, -7.565426e-20, -7.779635e-20, 2.9100894e-19, -9.0222664e-20, 4.4913103e-20, 2.2742708e-19, -9.628549e-20, 1.3589648e-19, 1.6628895e-19, -9.552959e-20, 1.976291e-19, 1.1042565e-19, -8.9620787e-20, 2.3362977e-19, 6.169972e-20, -8.011591e-20, 2.4801594e-19, 2.1131757e-20, -6.840185e-20, 2.4513117e-19, -1.0956079e-20, -5.565857e-20, 2.29249e-19, -3.479174e-20, -4.2842534e-20, 2.0435087e-19, -5.1009566e-20, -3.068651e-20, 1.7397356e-19, -6.051812e-20, -1.9711943e-20, 1.4111752e-19, -6.438416e-20, -1.02501645e-20, 1.08207134e-19, -6.373543e-20, -2.4691567e-21, 7.709257e-20, -5.9683175e-20, 3.5969246e-21, 4.9083156e-20, -5.326403e-20, 8.017791e-21, 2.5003132e-20, -4.539994e-20, 1.0938399e-20, 5.2611082e-21, -3.6873967e-20, 1.2552938e-20, -1.0073764e-20, -2.831968e-20, 1.30822726e-20, -2.1194828e-20, -2.0221351e-20, 1.27552535e-20, -2.848462e-20, -1.29225015e-20, 1.1794047e-20, -3.2448473e-20, -6.6402174e-21, 1.040332e-20, -3.3657058e-20, -1.4831455e-21, 8.762984e-21, -3.2698973e-20, 2.5287517e-21, 7.024046e-21, -3.0143618e-20, 5.4441942e-21, 5.307059e-21, -2.6513976e-20, 7.36151e-21, 3.702647e-21, -2.2268473e-20, 8.411334e-21, 2.2735693e-21, -1.7790757e-20, 8.741621e-21, 1.0578539e-21, -1.3386087e-20, 8.505266e-21, 7.256309e-23, -9.2829585e-21, 7.850388e-21, -6.8216713e-22, -5.6386253e-21, 6.9132016e-21, -1.219104e-21, -2.5472853e-21, 5.8132464e-21, -1.5601328e-21, -4.9835294e-23, 4.6506845e-21, -1.7328642e-21, 1.8557193e-21, 3.5053224e-21, -1.7677298e-21, 3.2039401e-21, 2.437004e-21, -1.6956106e-21, 4.0522726e-21, 1.4870224e-21, -1.5460074e-21, 4.472389e-21, 6.802325e-22, -1.3457218e-21, 4.5428012e-21, 2.757682e-23, -1.1180027e-21, 4.3428477e-21, -4.7121194e-22, -8.820947e-22, 3.948069e-21, -8.24927e-22, -6.5311725e-22, 3.426893e-21, -1.0483665e-21, -4.422025e-22, 2.8385119e-21, -1.1600774e-21, -2.5682378e-22, 2.2317739e-21, -1.1804276e-21, -1.0124925e-22, 1.6449211e-21, -1.1300353e-21, 2.2933018e-23, 1.1059793e-21, -1.0285586e-21, 1.1626554e-22, 6.336261e-22, -8.938261e-22, 1.8088382e-22, 2.3837498e-22, -7.412779e-22, 2.2001785e-22, -7.606852e-23, -5.83672e-22, 2.3755114e-22, -3.1139218e-22, -4.3101113e-22, 2.3764832e-22, -4.7329867e-22, -2.906399e-22, 2.244558e-22, -5.7023137e-22, -1.6746823e-22, 2.0187443e-22, -6.122501e-22, -6.4276595e-23, 1.7340047e-22, -6.100851e-22, 1.7931888e-23, 1.4202657e-22, -5.743779e-22, 7.9564347e-23, 1.1019467e-22, -5.151087e-22, 1.2207962e-22, 7.979081e-23, -4.4119665e-22, 1.4765638e-22, 5.2172263e-23, -3.602545e-22, 1.5890013e-22, 2.8217583e-23, -2.7847477e-22, 1.5859605e-22, 8.3916104e-24, -2.0062222e-22, 1.4951084e-22, -7.18198e-24, -1.3010781e-22, 1.3424258e-22, -1.8646351e-23, -6.912066e-23, 1.1511587e-22, -2.6339973e-23, -1.879677e-23, 9.4117215e-23, -3.0731222e-23, 2.0593626e-23, 7.286459e-23, -3.2361296e-23, 4.945499e-23, 5.2604874e-23, -3.1796676e-23, 6.8683266e-23, 3.4232638e-23, -2.9591466e-23, 7.949881e-23, 1.8324068e-23, -2.6259419e-23, 8.330104e-23, 5.1806176e-24, -2.2254858e-23, 8.1547676e-23, -5.1224004e-24, -1.7961473e-23, 7.565945e-23, -1.26861716e-23, -1.3687713e-23, 6.694964e-23, -1.7740704e-23, -9.667485e-24, 5.657633e-23, -2.0601317e-23, -6.064846e-24, 4.55147e-23, -2.1630719e-23, -2.9814785e-24, 3.4546163e-23, -2.1207483e-23, -4.6586417e-25, 2.4260867e-23, -1.9701127e-23, 1.4767541e-24, 1.507029e-23, -1.7453652e-23, 2.874369e-24, 7.226827e-24, -1.4766989e-23, 3.778732e-24, 8.475672e-25, -1.1895698e-23, 4.256808e-24, -4.0600174e-24, -9.044031e-24, 4.3834133e-24, -7.5723894e-24, -6.366506e-24, 4.23517e-24, -9.825692e-24, -3.97113e-24, 3.8857994e-24, -1.0993938e-23, -1.9244404e-24, 3.402696e-24, -1.1270277e-23, -2.5766485e-25, 2.8446725e-24, -1.0851658e-23, 1.0266122e-24, 2.2607198e-24, -9.92693e-24, 1.947775e-24, 1.6896105e-24, -8.668227e-24, 2.5408626e-24, 1.1601689e-24, -7.225339e-24, 2.8508855e-24, 6.9202867e-25, -5.7226715e-24, 2.9279383e-24, 2.9672705e-25, -4.258345e-24, 2.8231932e-24, -2.1012418e-26, -2.904975e-24, 2.5857859e-24, -2.619207e-25, -1.7116923e-24, 2.2605584e-24, -4.308438e-25, -7.069925e-25, 1.8865774e-24, -5.354923e-25, 9.794186e-26, 1.4963294e-24, -5.853289e-25, 7.057426e-25, 1.1154731e-24, -5.906231e-25, 1.12941985e-24, 7.630331e-25, -5.6168543e-25, 1.3891643e-24, 4.519181e-25, -5.082824e-25, 1.5095106e-24, 1.8965576e-25, -4.3922074e-25, 1.5169332e-24, -2.0745697e-26, -3.6208437e-25, 1.4379062e-24, -1.7988952e-25, -2.8310206e-25, 1.2974263e-24, -2.9109675e-25, -2.071225e-25, 1.1179684e-24, -3.5957367e-25, -1.3767223e-25, 9.18832e-25, -3.9167227e-25, -7.7073535e-26, 7.1581934e-25, -3.9426282e-25, -2.6601647e-26, 5.2118655e-25, -3.74227e-25, 1.3337208e-26, 3.4380358e-25, -3.3807098e-25, 4.3021525e-26, 1.8946527e-25, -2.9165154e-25, 6.323594e-26, 6.130027e-26, -2.4000393e-25, 7.5106904e-26, -3.9768928e-26, -1.8725623e-25, 7.9958424e-26, -1.1455207e-25, -1.36615e-25, 7.919109e-26, -1.6513349e-25, -9.040569e-26, 7.418566e-26, -1.9445228e-25, -5.0152606e-26, 6.623073e-26, -2.0593465e-25, -1.6684595e-26, 5.647267e-26, -2.0318672e-25, 9.745626e-27, 4.5885583e-26};
	localparam real hb[0:1199] = {0.09036497, 0.0042399773, -0.009115652, 0.085569896, 0.0101578925, -0.008072455, 0.07845638, 0.014705096, -0.0064387238, 0.06969149, 0.017824404, -0.004529465, 0.059936076, 0.019579753, -0.0025822371, 0.049796417, 0.02011784, -0.00076614704, 0.039793197, 0.019635536, 0.00080829044, 0.030344823, 0.018353287, 0.0020790123, 0.021762133, 0.016494296, 0.0030224824, 0.014251728, 0.014269142, 0.0036443763, 0.00792538, 0.0118652405, 0.0039711646, 0.0028133253, 0.009440502, 0.004042785, -0.0011204077, 0.0071204356, 0.0039065, -0.003962103, 0.004997996, 0.0036119597, -0.005833038, 0.003135466, 0.003207425, -0.0068755466, 0.0015677463, 0.002737062, -0.0072409683, 0.00030650996, 0.0022391828, -0.007079774, -0.0006552493, 0.0017452879, -0.0065339375, -0.0013386372, 0.0012797649, -0.0057314746, -0.0017745271, 0.00086008897, -0.004782968, -0.0019996704, 0.00049739145, -0.003779821, -0.0020533716, 0.00019726786, -0.0027939335, -0.001974784, -3.9279374e-05, -0.0018785027, -0.0018008389, -0.00021485309, -0.0010696395, -0.0015647728, -0.00033469673, -0.00038852476, -0.0012952005, -0.00040580356, 0.00015613581, -0.0010156557, -0.0004361338, 0.000565563, -0.0007445162, -0.000433959, 0.00084842165, -0.00049522973, -0.00040734102, 0.0010185246, -0.00027675464, -0.0003637436, 0.0010928051, -9.414373e-05, -0.00030976746, 0.0010896028, 5.0796905e-05, -0.00025099434, 0.0010272873, 0.00015882665, -0.00019192393, 0.0009232092, 0.0002326101, -0.00013598464, 0.0007929628, 0.00027610926, -8.560091e-05, 0.00064992433, 0.00029404912, -4.2299594e-05, 0.00050502596, 0.00029146875, -6.8407016e-06, 0.0003667219, 0.00027336265, 2.064079e-05, 0.00024110163, 0.00024441042, 4.049228e-05, 0.00013210971, 0.00020878887, 5.340824e-05, 4.1833468e-05, 0.0001700573, 6.030798e-05, -2.9173532e-05, 0.00013110481, 6.2230145e-05, -8.1558894e-05, 9.4147814e-05, 6.02458e-05, -0.00011685057, 6.0765855e-05, 5.5390527e-05, -0.00013716304, 3.196459e-05, 4.8614744e-05, -0.00014494038, 8.255933e-06, 4.0750678e-05, -0.0001427421, -1.02532995e-05, 3.2493856e-05, -0.00013307319, -2.3771094e-05, 2.4396679e-05, -0.00011825778, -3.273387e-05, 1.6871538e-05, -0.00010035267, -3.7727885e-05, 1.0201045e-05, -8.1096485e-05, -3.9420913e-05, 4.553076e-06, -6.188855e-05, -3.8505677e-05, -1.3351346e-09, -4.379175e-05, -3.5655296e-05, -3.4689465e-06, -2.7553384e-05, -3.149042e-05, -5.9154463e-06, -1.3638718e-05, -2.6557156e-05, -7.4477807e-06, -2.2722415e-06, -2.1314321e-05, -8.198382e-06, 6.5174827e-06, -1.6128675e-05, -8.311723e-06, 1.2852708e-05, -1.1276375e-05, -7.933403e-06, 1.6963733e-05, -6.9491484e-06, -7.201757e-06, 1.915029e-05, -3.2637115e-06, -6.241874e-06, 1.9748253e-05, -2.731218e-07, -5.1617753e-06, 1.910227e-05, 2.0210155e-06, -4.050452e-06, 1.7544417e-05, 3.6563804e-06, -2.977433e-06, 1.537864e-05, 4.6984746e-06, -1.9935424e-06, 1.2870485e-05, 5.2303367e-06, -1.1325161e-06, 1.0241401e-05, 5.343727e-06, -4.1319177e-07, 7.666878e-06, 5.131927e-06, 1.5799479e-07, 5.2775918e-06, 4.6841674e-06, 5.844146e-07, 3.16277e-06, 4.081608e-06, 8.767209e-07, 1.3750837e-06, 3.394731e-06, 1.0505199e-06, -6.359334e-08, 2.681946e-06, 1.1243196e-06, -1.1560729e-06, 1.9892025e-06, 1.1178051e-06, -1.9238194e-06, 1.3503931e-06, 1.0504591e-06, -2.4013098e-06, 7.883302e-07, 9.4052206e-07, -2.6310133e-06, 3.1611168e-07, 8.042696e-07, -2.6591165e-06, -6.129808e-08, 6.555715e-07, -2.5320603e-06, -3.454086e-07, 5.0569054e-07, -2.2938889e-06, -5.4257777e-07, 3.632738e-07, -1.9843594e-06, -6.625024e-07, 2.344932e-07, -1.6377461e-06, -7.168822e-07, 1.2328992e-07, -1.2822309e-06, -7.182897e-07, 3.1685722e-08, -9.3978184e-07, -6.7926067e-07, -3.9873004e-08, -6.264063e-07, -6.1160307e-07, -9.216509e-08, -3.5267666e-07, -5.259113e-07, -1.2685935e-07, -1.2443446e-07, -4.3126354e-07, -1.4620956e-07, 5.640928e-08, -3.3507646e-07, -1.5278935e-07, 1.910447e-07, -2.4308642e-07, -1.492724e-07, 2.8295824e-07, -1.5942956e-07, -1.3825932e-07, 3.3719118e-07, -8.679187e-08, -1.2214998e-07, 3.5968802e-07, -2.660465e-08, -1.0305723e-07, 3.567494e-07, 2.073672e-08, -8.275738e-08, 3.3459582e-07, 5.5648126e-08, -6.267113e-08, 2.9903916e-07, 7.914034e-08, -4.3868962e-08, 2.552557e-07, 9.2620944e-08, -2.7094774e-08, 2.076485e-07, 9.772125e-08, -1.28021105e-08, 1.5978559e-07, 9.615197e-08, -1.1979872e-09, 1.1439974e-07, 8.9588816e-08, 7.709966e-09, 7.3434734e-08, 7.958725e-08, 1.4066451e-08, 3.812472e-08, 6.752433e-08, 1.8124151e-08, 9.094313e-09, 5.4564296e-08, 2.020391e-08, -1.35311655e-08, 4.1644235e-08, 2.0660599e-08, -3.0013776e-08, 2.9475874e-08, 1.9855193e-08, -4.08961e-08, 1.8559513e-08, 1.8133171e-08, -4.690415e-08, 9.206431e-09, 1.5808924e-08, -4.8863175e-08, 1.5665158e-09, 1.3155593e-08, -4.7627942e-08, -4.3416697e-09, 1.039966e-08, -4.4028017e-08, -8.600654e-09, 7.719402e-09, -3.8827427e-08, -1.1365383e-08, 5.246423e-09, -3.2697635e-08, -1.283732e-08, 3.0694185e-09, -2.6202096e-08, -1.32421265e-08, 1.2394428e-09, -1.979051e-08, -1.2811306e-08, -2.239797e-10, -1.3800811e-08, -1.1767882e-08, -1.3264359e-09, -8.466915e-09, -1.0315974e-08, -2.0923332e-09, -3.9304298e-09, -8.633901e-09, -2.5590552e-09, -2.5472774e-10, -6.8703674e-09, -2.7717857e-09, 2.5599607e-09, -5.14322e-09, -2.7791278e-09, 4.5615254e-09, -3.5402123e-09, -2.6295779e-09, 5.8318466e-09, -2.1212718e-09, -2.3688427e-09, 6.4741275e-09, -9.2178154e-10, -2.0379525e-09, 6.602058e-09, 4.3551884e-11, -1.6720838e-09, 6.3309704e-09, 7.76595e-10, -1.2999902e-09, 5.77101e-09, 1.2917376e-09, -9.439258e-10, 5.0222204e-09, 1.6121071e-09, -6.19951e-10, 4.1713655e-09, 1.7661972e-09, -3.3851055e-10, 3.2902467e-09, 1.7849994e-09, -1.0518775e-10, 2.4352584e-09, 1.699678e-09, 7.844976e-11, 1.6479078e-09, 1.5397891e-09, 2.1398125e-10, 9.560427e-10, 1.332014e-09, 3.0529546e-10, 3.7554979e-10, 1.0993542e-09, 3.5782352e-10, -8.768451e-11, 8.60723e-10, 3.7786865e-10, -4.357213e-10, 6.308638e-10, 3.7204642e-10, -6.7656175e-10, 4.2051962e-10, 3.4684128e-10, -8.2228596e-10, 2.3678604e-10, 3.0827557e-10, -8.874075e-10, 8.3583536e-11, 2.616836e-10, -8.874836e-10, -3.7805332e-11, 2.1157745e-10, -8.379982e-10, -1.2817936e-10, 1.6159109e-10, -7.535152e-10, -1.898785e-10, 1.1448643e-10, -6.470841e-10, -2.2628636e-10, 7.220689e-11, -5.298726e-10, -2.4139268e-10, 3.5963798e-11, -4.1099088e-10, -2.3942634e-10, 6.343025e-12, -2.974732e-10, -2.2456235e-10, -1.6578725e-11, -1.9437936e-10, -2.0070161e-10, -3.311699e-11, -1.0498246e-10, -1.7131838e-10, -4.386852e-11, -3.101161e-11, -1.3936793e-10, -4.9611024e-11, 2.7076966e-11, -1.07245185e-10, -5.121665e-11, 6.982229e-11, -7.6784405e-11, -4.9580805e-11, 9.849156e-11, -4.9290304e-11, -4.5566658e-11, 1.1483604e-10, -2.5591326e-11, -3.9964598e-11, 1.2087802e-10, -6.106779e-12, -3.346546e-11, 1.1873334e-10, 9.079133e-12, -2.6645667e-11, 1.1047113e-10, 2.0142232e-11, -1.996228e-11, 9.800927e-11, 2.7446623e-11, -1.3755915e-11, 8.3043426e-11, 3.1479545e-11, -8.259455e-12, 6.7005304e-11, 3.279484e-11, -3.6106985e-12, 5.1045546e-11, 3.196619e-11, 1.3268992e-13, 3.6036434e-11, 2.955036e-11, 2.9773183e-12, 2.2589486e-11, 2.6060135e-11, 4.978394e-12, 1.1083396e-11, 2.1946188e-11, 6.2250695e-12, 1.6983405e-12, 1.7586694e-11, 6.827383e-12, -5.546812e-12, 1.3283488e-11, 6.905142e-12, -1.0757145e-11, 9.263391e-12, 6.578909e-12, -1.4126313e-11, 5.6834108e-12, 5.963093e-12, -1.590464e-11, 2.6386003e-12, 5.161024e-12, -1.6371656e-11, 1.7150272e-13, 4.2618274e-12, -1.581353e-11, -1.7177186e-12, 3.338828e-12, -1.4505517e-11, -3.0611995e-12, 2.449219e-12, -1.2699198e-11, -3.9138887e-12, 1.6347117e-12, -1.0614062e-11, -4.3450504e-12, 9.228931e-13, -8.432901e-12, -4.430986e-12, 3.2904823e-13, -6.3003426e-12, -4.2491015e-12, -1.4176282e-13, -4.3238624e-12, -3.8733222e-12, -4.9255337e-13, -2.576632e-12, -3.370795e-12, -7.323193e-13, -1.1016023e-12, -2.7997535e-12, -8.7411225e-13, 8.369866e-14, -2.2083902e-12, -9.333455e-13, 9.820906e-13, -1.6345563e-12, -9.263709e-13, 1.6117382e-12, -1.1061121e-12, -8.6934285e-13, 2.0014836e-12, -6.417495e-13, -7.7736336e-13, 2.1866933e-12, -2.5213284e-13, -6.6388957e-13, 2.205731e-12, 5.8785916e-14, -5.403741e-13, 2.0971016e-12, 2.923889e-13, -4.1610332e-13, 1.8972688e-12, 4.540453e-13, -2.9819436e-13, 1.639105e-12, 5.518622e-13, -1.9171462e-13, 1.3509112e-12, 5.955801e-13, -9.988681e-14, 1.0559265e-12, 5.9564024e-13, -2.434834e-14, 7.722352e-13, 5.6243476e-13, 3.4562603e-14, 5.1298505e-13, 5.0573825e-13, 7.751659e-14, 2.8682886e-13, 4.3430944e-13, 1.0591532e-13, 9.8511504e-14, 3.556437e-13, 1.2163924e-13, -5.0464227e-14, 2.7585573e-13, 1.2682863e-13, -1.6114962e-13, 1.9966689e-13, 1.2370221e-13, -2.364832e-13, 1.3047335e-13, 1.1441462e-13, -2.8067723e-13, 7.047216e-14, 1.0095139e-13, -2.986794e-13, 2.0824002e-14, 8.505839e-14, -2.9572137e-13, -1.8164727e-14, 6.8201385e-14, -2.769592e-13, -4.685566e-14, 5.1550964e-14, -2.4720344e-13, -6.609919e-14, 3.598743e-14, -2.1073295e-13, -7.707061e-14, 2.2120811e-14, -1.7118251e-13, -8.112716e-14, 1.0321143e-14, -1.3149341e-13, -7.968891e-14, 7.5496677e-16, -9.391428e-14, -7.414453e-14, -6.5755155e-15, -6.004055e-14, -6.5781256e-14, -1.1793434e-14, -3.088089e-14, -5.5737197e-14, -1.511053e-14, -6.9406384e-15, -4.4973262e-14, -1.6794243e-14, 1.1686564e-14, -3.426176e-14, -1.7139508e-14, 2.5225974e-14, -2.4188173e-14, -1.6445758e-14, 3.4133236e-14, -1.5162952e-14, -1.4999124e-14, 3.9014083e-14, -7.440298e-15, -1.3059634e-14, 4.0554792e-14, -1.1411637e-15, -1.0852915e-14, 3.9464685e-14, 3.721764e-15, -8.565789e-15, 3.6431053e-14, 7.218995e-15, -6.345079e-15, 3.2086025e-14, 9.480491e-15, -4.2989395e-15, 2.6984422e-14, 1.0674249e-14, -2.5000283e-15, 2.159119e-14, 1.0987872e-14, -9.898999e-16, 1.6276843e-14, 1.06134245e-14, 2.1590663e-16, 1.1319271e-14, 9.735649e-15, 1.122541e-15, 6.910272e-15, 8.523397e-15, 1.7506278e-15, 3.1653545e-15, 7.123984e-15, 2.1314305e-15, 1.3544979e-16, 5.660098e-15, 2.3025729e-15, -2.180554e-15, 4.2288116e-15, 2.3044236e-15, -3.823357e-15, 2.902263e-15, 2.1771906e-15, -4.8615486e-15, 1.7295667e-15, 1.9587129e-15, -5.381139e-15, 7.395535e-16, 1.6829136e-15, -5.476608e-15, -5.600905e-17, 1.3788382e-15, -5.243616e-15, -6.5901043e-16, 1.0701944e-15, -4.77338e-15, -1.0816399e-15, 7.752999e-16, -4.1486424e-15, -1.3432534e-15, 5.0734314e-16, -3.4410677e-15, -1.4675866e-15, 2.748684e-16, -2.7098803e-15, -1.4803871e-15, 8.240478e-17, -2.0015213e-15, -1.4074978e-15, -6.8830804e-17, -1.3500983e-15, -1.2733915e-15, -1.8021264e-16, -7.784197e-16, -1.1001314e-15, -2.5501264e-16, -2.994108e-16, -9.067127e-16, -2.9776578e-16, 8.2253894e-17, -7.087328e-16, -3.1371618e-16, 3.6844713e-16, -5.1833006e-16, -3.083555e-16, 5.659254e-16, -3.4432932e-16, -2.8705748e-16, 6.8478887e-16, -1.9253857e-16, -2.5480599e-16, 7.371213e-16, -6.614294e-17, -2.160096e-16, 7.358432e-16, 3.3848535e-17, -1.7439256e-16, 6.937914e-16, 1.08141074e-16, -1.3294972e-16, 6.230221e-16, 1.587066e-16, -9.395315e-17, 5.343241e-16, 1.8837207e-16, -5.899732e-17, 4.3691796e-16, 2.0045798e-16, -2.907146e-17, 3.3831483e-16, 1.9847562e-16, -4.6484643e-18, 2.443042e-16, 1.8588548e-16, 1.4218575e-17, 1.5904068e-16, 1.6591627e-16, 2.7799367e-17, 8.520121e-17, 1.414398e-16, 3.6594497e-17, 2.4187628e-17, 1.1489572e-16, 4.1252513e-17, -2.3648035e-17, 8.825816e-17, 4.2498492e-17, -5.877322e-17, 6.3036404e-17, 4.107533e-17, -8.225363e-17, 4.030132e-17, 3.7698032e-17, -9.555126e-17, 2.0729977e-17, 3.302044e-17, -1.00348437e-16, 4.6616007e-18, 2.76133e-17, -9.840144e-17, -7.840903e-18, 2.1952177e-17, -9.142484e-17, -1.6928673e-17, 1.6413576e-17, -8.100571e-17, -2.2907483e-17, 1.1277513e-17, -6.8545427e-17, -2.6183858e-17, 6.7348566e-18, -5.5225592e-17, -2.7218381e-17, 2.8978999e-18, -4.1994454e-17, -2.6487117e-17, -1.8719799e-19, -2.9569517e-17, -2.4451348e-17, -2.527241e-18, -1.8452424e-17, -2.153534e-17, -4.169005e-18, -8.952369e-18, -1.8111474e-17, -5.1871102e-18, -1.2146473e-18, -1.4491814e-17, -5.6732224e-18, 4.7484224e-18, -1.0925047e-17, -5.7268795e-18, 9.026524e-18, -7.597691e-18, -5.44806e-18, 1.178205e-17, -4.638488e-18, -4.931496e-18, 1.3223719e-17, -2.124971e-18, -4.262635e-18, 1.3583899e-17, -9.133178e-20, -3.5150796e-18, 1.31000015e-17, 1.4631681e-18, -2.7493e-18, 1.2000025e-17, 2.5658394e-18, -2.0123846e-18, 1.0492073e-17, 3.2627128e-18, -1.3385989e-18, 8.757471e-18, 3.6115115e-18, -7.5052423e-19, 6.94702e-18, 3.6756457e-18, -2.6058066e-19, 5.179849e-18, 3.5193173e-18, 1.2724733e-19, 3.544303e-18, 3.203749e-18, 4.1562455e-19, 2.1003448e-18, 2.7844742e-18, 6.1213314e-19, 8.829621e-19, 2.3095925e-18, 7.276783e-19, -9.3835756e-20, 1.818855e-18, 7.7508824e-19, -8.328061e-19, 1.3434323e-18, 7.679403e-19, -1.3493264e-18, 9.062178e-19, 7.1962454e-19, -1.6675306e-18, 5.225211e-19, 6.426407e-19, -1.8168768e-18, 2.0101838e-19, 5.481127e-19, -1.8292355e-18, -5.5151815e-20, 4.45495e-19, -1.7365352e-18, -2.4724553e-19, 3.4244254e-19, -1.5689669e-18, -3.7979667e-19, 2.4481157e-19, -1.3537122e-18, -4.595836e-19, 1.567614e-19, -1.1141423e-18, -4.9471615e-19, 8.0926084e-20, -8.694209e-19, -4.9386586e-19, 1.8630547e-20, -6.3443605e-19, -4.656482e-19, -2.98716e-20, -4.199873e-19, -4.18155e-19, -6.515714e-20, -2.331562e-19, -3.586273e-19, -8.840334e-20, -7.779635e-20, -2.9325378e-19, -1.0117923e-19, 4.4913103e-20, -2.2707586e-19, -1.0526472e-19, 1.3589648e-19, -1.6397942e-19, -1.0250104e-19, 1.976291e-19, -1.06753054e-19, -9.4673374e-20, 2.3362977e-19, -5.719364e-20, -8.3424486e-20, 2.4801594e-19, -1.624221e-20, -7.019698e-20, 2.4513117e-19, 1.5864831e-20, -5.620042e-20, 2.29249e-19, 3.9441093e-20, -4.2399275e-20, 2.0435087e-19, 5.520174e-20, -2.9517455e-20, 1.7397356e-19, 6.412795e-20, -1.805518e-20, 1.4111752e-19, 6.7348793e-20, -8.314308e-21, 1.08207134e-19, 6.6043e-20, -4.287322e-22, 7.709257e-20, 6.136131e-20, 5.6031127e-21, 4.9083156e-20, 5.436894e-20, 9.8859005e-21, 2.5003132e-20, 4.6006425e-20, 1.2597021e-20, 5.2611082e-21, 3.7066858e-20, 1.3959364e-20, -1.0073764e-20, 2.8186687e-20, 1.4218041e-20, -2.1194828e-20, 1.98475e-20, 1.3621408e-20, -2.848462e-20, 1.2386013e-20, 1.2406432e-20, -3.2448473e-20, 6.009766e-21, 1.0788177e-20, -3.3657058e-20, 8.1630034e-22, 8.9530055e-21, -3.2698973e-20, -3.1860986e-21, 7.055018e-21, -3.0143618e-20, -6.0576084e-21, 5.2151238e-21, -2.6513976e-20, -7.907209e-21, 3.522203e-21, -2.2268473e-20, -8.874978e-21, 2.0357644e-21, -1.7790757e-20, -9.1168664e-21, 7.8962225e-22, -1.3386087e-20, -8.792213e-21, -2.0387647e-22, -9.2829585e-21, -8.054044e-21, -9.494281e-22, -5.6386253e-21, -7.04203e-21, -1.4644521e-21, -2.5472853e-21, -5.8778727e-21, -1.7750894e-21, -4.9835294e-23, -4.6627884e-21, -1.9126663e-21, 1.8557193e-21, -3.4767346e-21, -1.9107105e-21, 3.2039401e-21, -2.3790096e-21, -1.802556e-21, 4.0522726e-21, -1.4098612e-21, -1.6195278e-21, 4.472389e-21, -5.927757e-22, -1.3896718e-21, 4.5428012e-21, 6.284181e-23, -1.13697e-21, 4.3428477e-21, 5.5883957e-22, -8.809692e-22, 3.948069e-21, 9.055364e-22, -6.367461e-22, 3.426893e-21, 1.1191288e-21, -4.1512989e-22, 2.8385119e-21, 1.2193871e-21, -2.2310915e-22, 2.2317739e-21, 1.2277008e-21, -6.435626e-23, 1.6449211e-21, 1.1654992e-21, 6.018802e-23, 1.1059793e-21, 1.0530451e-21, 1.5171661e-22, 6.336261e-22, 9.085823e-22, 2.1298146e-22, 2.3837498e-22, 7.477969e-22, 2.4776871e-22, -7.606852e-23, 5.835514e-22, 2.604411e-22, -3.1139218e-22, 4.258385e-22, 2.55557e-22, -4.7329867e-22, 2.8190703e-22, 2.3756954e-22, -5.7023137e-22, 1.5651034e-22, 2.1060294e-22, -6.122501e-22, 5.223523e-23, 1.7830065e-22, -6.100851e-22, -3.0126538e-23, 1.4373645e-22, -5.743779e-22, -9.119503e-23, 1.0937845e-22, -5.151087e-22, -1.3263135e-22, 7.709557e-23, -4.4119665e-22, -1.5679702e-22, 4.8195867e-23, -3.602545e-22, -1.664554e-22, 2.3487078e-23, -2.7847477e-22, -1.6452169e-22, 3.3506394e-24, -2.0062222e-22, -1.5386409e-22, -1.2178081e-23, -1.3010781e-22, -1.3715483e-22, -2.3329362e-23, -6.912066e-23, -1.1676767e-22, -3.052302e-23, -1.879677e-23, -9.471648e-23, -3.4299833e-23, 2.0593626e-23, -7.2628486e-23, -3.5262565e-23, 4.945499e-23, -5.17455e-23, -3.4027544e-23, 6.8683266e-23, -3.2946378e-23, -3.1187026e-23, 7.949881e-23, -1.6784373e-23, -2.7281874e-23, 8.330104e-23, -3.5337864e-24, -2.2783597e-23, 8.1547676e-23, 6.758923e-24, -1.808454e-23, 7.565945e-23, 1.4223482e-23, -1.3494832e-23, 6.694964e-23, 1.9116607e-23, -9.244656e-24, 5.657633e-23, 2.1777436e-23, -5.4904273e-24, 4.55147e-23, 2.258897e-23, -2.3236324e-24, 3.4546163e-23, 2.194625e-23, 2.188204e-25, 2.4260867e-23, 2.0231431e-23, 2.1436642e-24, 1.507029e-23, 1.7795525e-23, 3.490507e-24, 7.226827e-24, 1.4946215e-23, 4.3217922e-24, 8.475672e-25, 1.1941002e-23, 4.713875e-24, -4.0600174e-24, 8.98477e-24, 4.7494475e-24, -7.5723894e-24, 6.230888e-24, 4.5114143e-24, -9.825692e-24, 3.7849077e-24, 4.0782125e-24, -1.0993938e-23, 1.7100586e-24, 3.520498e-24, -1.1270277e-23, 3.3796607e-26, 2.8990532e-24, -1.0851658e-23, -1.2452107e-24, 2.2637446e-24, -9.92693e-24, -2.1501554e-24, 1.65333965e-24, -8.668227e-24, -2.7195889e-24, 1.0959836e-24, -7.225339e-24, -3.0016126e-24, 6.10159e-25, -5.7226715e-24, -3.048919e-24, 2.059542e-25, -4.258345e-24, -2.9147568e-24, -1.1350111e-25, -2.904975e-24, -2.6498256e-24, -3.5055354e-25, -1.7116923e-24, -2.3000531e-24, -5.11591e-25, -7.069925e-25, -1.905167e-24, -6.0572394e-25, 9.794186e-26, -1.4979536e-24, -6.4362826e-25, 7.057426e-25, -1.1040809e-24, -6.365768e-25, 1.12941985e-24, -7.423601e-25, -5.956678e-25, 1.3891643e-24, -4.253281e-25, -5.31247e-25, 1.5095106e-24, -1.6004212e-25, -4.5250905e-25, 1.5169332e-24, 5.100987e-26, -3.672586e-25, 1.4379062e-24, 2.0895984e-25, -2.8180545e-25, 1.2974263e-24, 3.1763467e-25, -2.0096824e-25, 1.1179684e-24, 3.827007e-25, -1.2816054e-25, 9.18832e-25, 4.1090954e-25, -6.5534866e-26, 7.1581934e-25, 4.0946264e-25, -1.4162782e-26, 5.2118655e-25, 3.8550222e-25, 2.5767525e-26, 3.4380358e-25, 3.4572665e-25, 5.475141e-26, 1.8946527e-25, 2.9612216e-25, 7.377736e-26, 6.130027e-26, 2.4179834e-25, 8.415439e-26, -3.9768928e-26, 1.869115e-25, 8.7362617e-26, -1.1455207e-25, 1.3465973e-25, 8.4929955e-26, -1.6513349e-25, 8.733252e-26, 7.833537e-26, -1.9445228e-25, 4.6399285e-26, 6.893801e-26, -2.0593465e-25, 1.2622606e-26, 5.7929865e-26, -2.0318672e-25, -1.3816028e-26, 4.6309007e-26};
endpackage
